// this module implements a combo of sbox and tbox for a whole column
module direct_sbox_tbox(in_word, out_words);

input [0:31] in_word;
output [0:79] out_words[0:3];

wire [0:79] sbox_tbox[0:255];
wire [7:0] in_byte[0:3];
wire [0:79] mapping[0:3];

genvar i;
generate
    for(i = 0; i < 4; i++)
        begin: split_and_mapping
        // split original 32-bit column word into 4 bytes
        assign in_byte[i] = in_word[i*8:(i+1)*8-1];
        // map the "addresses" to the correct rom entry
        assign mapping[i] = sbox_tbox[in_byte[i]];
        end
endgenerate

assign out_words[0] = mapping[0];
assign out_words[1] = {mapping[1][0:7], mapping[1][8:39] >> 8 | mapping[1][8:39] << 24, mapping[1][40:47], mapping[1][48:79] >> 8 | mapping[1][48:79] << 24};
assign out_words[2] = {mapping[2][0:7], mapping[2][8:39] >> 16 | mapping[2][8:39] << 16, mapping[2][40:47], mapping[2][48:79] >> 16 | mapping[2][48:79] << 16};
assign out_words[3] = {mapping[3][0:7], mapping[3][8:39] >> 24 | mapping[3][8:39] << 8, mapping[3][40:47], mapping[3][48:79] >> 24 | mapping[3][48:79] << 8};

// hardwired implementation of the sbox_tbox mapping
assign sbox_tbox[0] = 80'h63c66363a55251f4a750;
assign sbox_tbox[1] = 80'h7cf87c7c84097e416553;
assign sbox_tbox[2] = 80'h77ee7777996a1a17a4c3;
assign sbox_tbox[3] = 80'h7bf67b7b8dd53a275e96;
assign sbox_tbox[4] = 80'hf2fff2f20d303bab6bcb;
assign sbox_tbox[5] = 80'h6bd66b6bbd361f9d45f1;
assign sbox_tbox[6] = 80'h6fde6f6fb1a5acfa58ab;
assign sbox_tbox[7] = 80'hc591c5c554384be30393;
assign sbox_tbox[8] = 80'h3060303050bf2030fa55;
assign sbox_tbox[9] = 80'h010201010340ad766df6;
assign sbox_tbox[10] = 80'h67ce6767a9a388cc7691;
assign sbox_tbox[11] = 80'h2b562b2b7d9ef5024c25;
assign sbox_tbox[12] = 80'hfee7fefe19814fe5d7fc;
assign sbox_tbox[13] = 80'hd7b5d7d762f3c52acbd7;
assign sbox_tbox[14] = 80'hab4dababe6d726354480;
assign sbox_tbox[15] = 80'h76ec76769afbb562a38f;
assign sbox_tbox[16] = 80'hca8fcaca457cdeb15a49;
assign sbox_tbox[17] = 80'h821f82829de325ba1b67;
assign sbox_tbox[18] = 80'hc989c9c9403945ea0e98;
assign sbox_tbox[19] = 80'h7dfa7d7d87825dfec0e1;
assign sbox_tbox[20] = 80'hfaeffafa159bc32f7502;
assign sbox_tbox[21] = 80'h59b25959eb2f814cf012;
assign sbox_tbox[22] = 80'h478e4747c9ff8d4697a3;
assign sbox_tbox[23] = 80'hf0fbf0f00b876bd3f9c6;
assign sbox_tbox[24] = 80'had41adadec34038f5fe7;
assign sbox_tbox[25] = 80'hd4b3d4d4678e15929c95;
assign sbox_tbox[26] = 80'ha25fa2a2fd43bf6d7aeb;
assign sbox_tbox[27] = 80'haf45afafea44955259da;
assign sbox_tbox[28] = 80'h9c239c9cbfc4d4be832d;
assign sbox_tbox[29] = 80'ha453a4a4f7de587421d3;
assign sbox_tbox[30] = 80'h72e4727296e949e06929;
assign sbox_tbox[31] = 80'hc09bc0c05bcb8ec9c844;
assign sbox_tbox[32] = 80'hb775b7b7c25475c2896a;
assign sbox_tbox[33] = 80'hfde1fdfd1c7bf48e7978;
assign sbox_tbox[34] = 80'h933d9393ae9499583e6b;
assign sbox_tbox[35] = 80'h264c26266a3227b971dd;
assign sbox_tbox[36] = 80'h366c36365aa6bee14fb6;
assign sbox_tbox[37] = 80'h3f7e3f3f41c2f088ad17;
assign sbox_tbox[38] = 80'hf7f5f7f70223c920ac66;
assign sbox_tbox[39] = 80'hcc83cccc4f3d7dce3ab4;
assign sbox_tbox[40] = 80'h346834345cee63df4a18;
assign sbox_tbox[41] = 80'ha551a5a5f44ce51a3182;
assign sbox_tbox[42] = 80'he5d1e5e5349597513360;
assign sbox_tbox[43] = 80'hf1f9f1f1080b62537f45;
assign sbox_tbox[44] = 80'h71e271719342b16477e0;
assign sbox_tbox[45] = 80'hd8abd8d873fabb6bae84;
assign sbox_tbox[46] = 80'h3162313153c3fe81a01c;
assign sbox_tbox[47] = 80'h152a15153f4ef9082b94;
assign sbox_tbox[48] = 80'h040804040c0870486858;
assign sbox_tbox[49] = 80'hc795c7c7522e8f45fd19;
assign sbox_tbox[50] = 80'h2346232365a194de6c87;
assign sbox_tbox[51] = 80'hc39dc3c35e66527bf8b7;
assign sbox_tbox[52] = 80'h183018182828ab73d323;
assign sbox_tbox[53] = 80'h96379696a1d9724b02e2;
assign sbox_tbox[54] = 80'h050a05050f24e31f8f57;
assign sbox_tbox[55] = 80'h9a2f9a9ab5b26655ab2a;
assign sbox_tbox[56] = 80'h070e07070976b2eb2807;
assign sbox_tbox[57] = 80'h12241212365b2fb5c203;
assign sbox_tbox[58] = 80'h801b80809ba286c57b9a;
assign sbox_tbox[59] = 80'he2dfe2e23d49d33708a5;
assign sbox_tbox[60] = 80'hebcdebeb266d302887f2;
assign sbox_tbox[61] = 80'h274e2727698b23bfa5b2;
assign sbox_tbox[62] = 80'hb27fb2b2cdd102036aba;
assign sbox_tbox[63] = 80'h75ea75759f25ed16825c;
assign sbox_tbox[64] = 80'h091209091b728acf1c2b;
assign sbox_tbox[65] = 80'h831d83839ef8a779b492;
assign sbox_tbox[66] = 80'h2c582c2c74f6f307f2f0;
assign sbox_tbox[67] = 80'h1a341a1a2e644e69e2a1;
assign sbox_tbox[68] = 80'h1b361b1b2d8665daf4cd;
assign sbox_tbox[69] = 80'h6edc6e6eb2680605bed5;
assign sbox_tbox[70] = 80'h5ab45a5aee98d134621f;
assign sbox_tbox[71] = 80'ha05ba0a0fb16c4a6fe8a;
assign sbox_tbox[72] = 80'h52a45252f6d4342e539d;
assign sbox_tbox[73] = 80'h3b763b3b4da4a2f355a0;
assign sbox_tbox[74] = 80'hd6b7d6d6615c058ae132;
assign sbox_tbox[75] = 80'hb37db3b3cecca4f6eb75;
assign sbox_tbox[76] = 80'h295229297b5d0b83ec39;
assign sbox_tbox[77] = 80'he3dde3e33e654060efaa;
assign sbox_tbox[78] = 80'h2f5e2f2f71b65e719f06;
assign sbox_tbox[79] = 80'h841384849792bd6e1051;
assign sbox_tbox[80] = 80'h53a65353f56c3e218af9;
assign sbox_tbox[81] = 80'hd1b9d1d1687096dd063d;
assign sbox_tbox[82] = 80'h000000000048dd3e05ae;
assign sbox_tbox[83] = 80'hedc1eded2c504de6bd46;
assign sbox_tbox[84] = 80'h2040202060fd91548db5;
assign sbox_tbox[85] = 80'hfce3fcfc1fed71c45d05;
assign sbox_tbox[86] = 80'hb179b1b1c8b90406d46f;
assign sbox_tbox[87] = 80'h5bb65b5bedda605015ff;
assign sbox_tbox[88] = 80'h6ad46a6abe5e1998fb24;
assign sbox_tbox[89] = 80'hcb8dcbcb4615d6bde997;
assign sbox_tbox[90] = 80'hbe67bebed946894043cc;
assign sbox_tbox[91] = 80'h397239394b5767d99e77;
assign sbox_tbox[92] = 80'h4a944a4adea7b0e842bd;
assign sbox_tbox[93] = 80'h4c984c4cd48d07898b88;
assign sbox_tbox[94] = 80'h58b05858e89de7195b38;
assign sbox_tbox[95] = 80'hcf85cfcf4a8479c8eedb;
assign sbox_tbox[96] = 80'hd0bbd0d06b90a17c0a47;
assign sbox_tbox[97] = 80'hefc5efef2ad87c420fe9;
assign sbox_tbox[98] = 80'haa4faaaae5abf8841ec9;
assign sbox_tbox[99] = 80'hfbedfbfb160000000000;
assign sbox_tbox[100] = 80'h43864343c58c09808683;
assign sbox_tbox[101] = 80'h4d9a4d4dd7bc322bed48;
assign sbox_tbox[102] = 80'h3366333355d31e1170ac;
assign sbox_tbox[103] = 80'h85118585940a6c5a724e;
assign sbox_tbox[104] = 80'h458a4545cff7fd0efffb;
assign sbox_tbox[105] = 80'hf9e9f9f910e40f853856;
assign sbox_tbox[106] = 80'h0204020206583daed51e;
assign sbox_tbox[107] = 80'h7ffe7f7f8105362d3927;
assign sbox_tbox[108] = 80'h50a05050f0b80a0fd964;
assign sbox_tbox[109] = 80'h3c783c3c44b3685ca621;
assign sbox_tbox[110] = 80'h9f259f9fba459b5b54d1;
assign sbox_tbox[111] = 80'ha84ba8a8e30624362e3a;
assign sbox_tbox[112] = 80'h51a25151f3d00c0a67b1;
assign sbox_tbox[113] = 80'ha35da3a3fe2c9357e70f;
assign sbox_tbox[114] = 80'h40804040c01eb4ee96d2;
assign sbox_tbox[115] = 80'h8f058f8f8a8f1b9b919e;
assign sbox_tbox[116] = 80'h923f9292adca80c0c54f;
assign sbox_tbox[117] = 80'h9d219d9dbc3f61dc20a2;
assign sbox_tbox[118] = 80'h38703838480f5a774b69;
assign sbox_tbox[119] = 80'hf5f1f5f504021c121a16;
assign sbox_tbox[120] = 80'hbc63bcbcdfc1e293ba0a;
assign sbox_tbox[121] = 80'hb677b6b6c1afc0a02ae5;
assign sbox_tbox[122] = 80'hdaafdada75bd3c22e043;
assign sbox_tbox[123] = 80'h214221216303121b171d;
assign sbox_tbox[124] = 80'h1020101030010e090d0b;
assign sbox_tbox[125] = 80'hffe5ffff1a13f28bc7ad;
assign sbox_tbox[126] = 80'hf3fdf3f30e8a2db6a8b9;
assign sbox_tbox[127] = 80'hd2bfd2d26d6b141ea9c8;
assign sbox_tbox[128] = 80'hcd81cdcd4c3a57f11985;
assign sbox_tbox[129] = 80'h0c180c0c1491af75074c;
assign sbox_tbox[130] = 80'h132613133511ee99ddbb;
assign sbox_tbox[131] = 80'hecc3ecec2f41a37f60fd;
assign sbox_tbox[132] = 80'h5fbe5f5fe14ff701269f;
assign sbox_tbox[133] = 80'h97359797a2675c72f5bc;
assign sbox_tbox[134] = 80'h44884444ccdc44663bc5;
assign sbox_tbox[135] = 80'h172e171739ea5bfb7e34;
assign sbox_tbox[136] = 80'hc493c4c457978b432976;
assign sbox_tbox[137] = 80'ha755a7a7f2f2cb23c6dc;
assign sbox_tbox[138] = 80'h7efc7e7e82cfb6edfc68;
assign sbox_tbox[139] = 80'h3d7a3d3d47ceb8e4f163;
assign sbox_tbox[140] = 80'h64c86464acf0d731dcca;
assign sbox_tbox[141] = 80'h5dba5d5de7b442638510;
assign sbox_tbox[142] = 80'h193219192be613972240;
assign sbox_tbox[143] = 80'h73e67373957384c61120;
assign sbox_tbox[144] = 80'h60c06060a096854a247d;
assign sbox_tbox[145] = 80'h8119818198acd2bb3df8;
assign sbox_tbox[146] = 80'h4f9e4f4fd174aef93211;
assign sbox_tbox[147] = 80'hdca3dcdc7f22c729a16d;
assign sbox_tbox[148] = 80'h2244222266e71d9e2f4b;
assign sbox_tbox[149] = 80'h2a542a2a7eaddcb230f3;
assign sbox_tbox[150] = 80'h903b9090ab350d8652ec;
assign sbox_tbox[151] = 80'h880b8888838577c1e3d0;
assign sbox_tbox[152] = 80'h468c4646cae22bb3166c;
assign sbox_tbox[153] = 80'heec7eeee29f9a970b999;
assign sbox_tbox[154] = 80'hb86bb8b8d337119448fa;
assign sbox_tbox[155] = 80'h142814143ce847e96422;
assign sbox_tbox[156] = 80'hdea7dede791ca8fc8cc4;
assign sbox_tbox[157] = 80'h5ebc5e5ee275a0f03f1a;
assign sbox_tbox[158] = 80'h0b160b0b1ddf567d2cd8;
assign sbox_tbox[159] = 80'hdbaddbdb766e223390ef;
assign sbox_tbox[160] = 80'he0dbe0e03b4787494ec7;
assign sbox_tbox[161] = 80'h3264323256f1d938d1c1;
assign sbox_tbox[162] = 80'h3a743a3a4e1a8ccaa2fe;
assign sbox_tbox[163] = 80'h0a140a0a1e7198d40b36;
assign sbox_tbox[164] = 80'h49924949db1da6f581cf;
assign sbox_tbox[165] = 80'h060c06060a29a57ade28;
assign sbox_tbox[166] = 80'h244824246cc5dab78e26;
assign sbox_tbox[167] = 80'h5cb85c5ce4893fadbfa4;
assign sbox_tbox[168] = 80'hc29fc2c25d6f2c3a9de4;
assign sbox_tbox[169] = 80'hd3bdd3d36eb75078920d;
assign sbox_tbox[170] = 80'hac43acacef626a5fcc9b;
assign sbox_tbox[171] = 80'h62c46262a60e547e4662;
assign sbox_tbox[172] = 80'h91399191a8aaf68d13c2;
assign sbox_tbox[173] = 80'h95319595a41890d8b8e8;
assign sbox_tbox[174] = 80'he4d3e4e437be2e39f75e;
assign sbox_tbox[175] = 80'h79f279798b1b82c3aff5;
assign sbox_tbox[176] = 80'he7d5e7e732fc9f5d80be;
assign sbox_tbox[177] = 80'hc88bc8c8435669d0937c;
assign sbox_tbox[178] = 80'h376e3737593e6fd52da9;
assign sbox_tbox[179] = 80'h6dda6d6db74bcf2512b3;
assign sbox_tbox[180] = 80'h8d018d8d8cc6c8ac993b;
assign sbox_tbox[181] = 80'hd5b1d5d564d210187da7;
assign sbox_tbox[182] = 80'h4e9c4e4ed279e89c636e;
assign sbox_tbox[183] = 80'ha949a9a9e020db3bbb7b;
assign sbox_tbox[184] = 80'h6cd86c6cb49acd267809;
assign sbox_tbox[185] = 80'h56ac5656fadb6e5918f4;
assign sbox_tbox[186] = 80'hf4f3f4f407c0ec9ab701;
assign sbox_tbox[187] = 80'heacfeaea25fe834f9aa8;
assign sbox_tbox[188] = 80'h65ca6565af78e6956e65;
assign sbox_tbox[189] = 80'h7af47a7a8ecdaaffe67e;
assign sbox_tbox[190] = 80'hae47aeaee95a21bccf08;
assign sbox_tbox[191] = 80'h0810080818f4ef15e8e6;
assign sbox_tbox[192] = 80'hba6fbabad51fbae79bd9;
assign sbox_tbox[193] = 80'h78f0787888dd4a6f36ce;
assign sbox_tbox[194] = 80'h254a25256fa8ea9f09d4;
assign sbox_tbox[195] = 80'h2e5c2e2e723329b07cd6;
assign sbox_tbox[196] = 80'h1c381c1c248831a4b2af;
assign sbox_tbox[197] = 80'ha657a6a6f1072a3f2331;
assign sbox_tbox[198] = 80'hb473b4b4c7c7c6a59430;
assign sbox_tbox[199] = 80'hc697c6c6513135a266c0;
assign sbox_tbox[200] = 80'he8cbe8e823b1744ebc37;
assign sbox_tbox[201] = 80'hdda1dddd7c12fc82caa6;
assign sbox_tbox[202] = 80'h74e874749c10e090d0b0;
assign sbox_tbox[203] = 80'h1f3e1f1f215933a7d815;
assign sbox_tbox[204] = 80'h4b964b4bdd27f104984a;
assign sbox_tbox[205] = 80'hbd61bdbddc8041ecdaf7;
assign sbox_tbox[206] = 80'h8b0d8b8b86ec7fcd500e;
assign sbox_tbox[207] = 80'h8a0f8a8a855f1791f62f;
assign sbox_tbox[208] = 80'h70e070709060764dd68d;
assign sbox_tbox[209] = 80'h3e7c3e3e425143efb04d;
assign sbox_tbox[210] = 80'hb571b5b5c47fccaa4d54;
assign sbox_tbox[211] = 80'h66cc6666aaa9e49604df;
assign sbox_tbox[212] = 80'h48904848d8199ed1b5e3;
assign sbox_tbox[213] = 80'h0306030305b54c6a881b;
assign sbox_tbox[214] = 80'hf6f7f6f6014ac12c1fb8;
assign sbox_tbox[215] = 80'h0e1c0e0e120d4665517f;
assign sbox_tbox[216] = 80'h61c26161a32d9d5eea04;
assign sbox_tbox[217] = 80'h356a35355fe5018c355d;
assign sbox_tbox[218] = 80'h57ae5757f97afa877473;
assign sbox_tbox[219] = 80'hb969b9b9d09ffb0b412e;
assign sbox_tbox[220] = 80'h861786869193b3671d5a;
assign sbox_tbox[221] = 80'hc199c1c158c992dbd252;
assign sbox_tbox[222] = 80'h1d3a1d1d279ce9105633;
assign sbox_tbox[223] = 80'h9e279e9eb9ef6dd64713;
assign sbox_tbox[224] = 80'he1d9e1e138a09ad7618c;
assign sbox_tbox[225] = 80'hf8ebf8f813e037a10c7a;
assign sbox_tbox[226] = 80'h982b9898b33b59f8148e;
assign sbox_tbox[227] = 80'h11221111334deb133c89;
assign sbox_tbox[228] = 80'h69d26969bbaecea927ee;
assign sbox_tbox[229] = 80'hd9a9d9d9702ab761c935;
assign sbox_tbox[230] = 80'h8e078e8e89f5e11ce5ed;
assign sbox_tbox[231] = 80'h94339494a7b07a47b13c;
assign sbox_tbox[232] = 80'h9b2d9b9bb6c89cd2df59;
assign sbox_tbox[233] = 80'h1e3c1e1e22eb55f2733f;
assign sbox_tbox[234] = 80'h8715878792bb1814ce79;
assign sbox_tbox[235] = 80'he9c9e9e9203c73c737bf;
assign sbox_tbox[236] = 80'hce87cece498353f7cdea;
assign sbox_tbox[237] = 80'h55aa5555ff535ffdaa5b;
assign sbox_tbox[238] = 80'h285028287899df3d6f14;
assign sbox_tbox[239] = 80'hdfa5dfdf7a617844db86;
assign sbox_tbox[240] = 80'h8c038c8c8f17caaff381;
assign sbox_tbox[241] = 80'ha159a1a1f82bb968c43e;
assign sbox_tbox[242] = 80'h8909898980043824342c;
assign sbox_tbox[243] = 80'h0d1a0d0d177ec2a3405f;
assign sbox_tbox[244] = 80'hbf65bfbfdaba161dc372;
assign sbox_tbox[245] = 80'he6d7e6e63177bce2250c;
assign sbox_tbox[246] = 80'h42844242c6d6283c498b;
assign sbox_tbox[247] = 80'h68d06868b826ff0d9541;
assign sbox_tbox[248] = 80'h41824141c3e139a80171;
assign sbox_tbox[249] = 80'h99299999b069080cb3de;
assign sbox_tbox[250] = 80'h2d5a2d2d7714d8b4e49c;
assign sbox_tbox[251] = 80'h0f1e0f0f11636456c190;
assign sbox_tbox[252] = 80'hb07bb0b0cb557bcb8461;
assign sbox_tbox[253] = 80'h54a85454fc21d532b670;
assign sbox_tbox[254] = 80'hbb6dbbbbd60c486c5c74;
assign sbox_tbox[255] = 80'h162c16163a7dd0b85742;

endmodule