module hardwired_sbox(in_word, out_word);

input [31:0] in_word;
output [31:0] out_word;

wire [7:0] sbox[255:0];
wire [7:0] in_byte[3:0];
wire [7:0] mapping[3:0];

genvar i;
generate
    for(i = 0; i < 4; i++)
        begin: packing_and_unpacking_words
        // unpack the input 32-bit word in 8-bit parts
        assign in_byte[i] = in_word[8*(i+1)-1:8*i];
        // pack the results of the sbox into a 32-bit word
        assign out_word[8*(i+1)-1:8*i] = mapping[i];
        // map in_addr to the output of sboxes
        assign mapping[i] = sbox[in_byte[i]];
        end
endgenerate

// hardwired implementation of the sbox
assign sbox[0] = 8'h63;
assign sbox[1] = 8'h7c;
assign sbox[2] = 8'h77;
assign sbox[3] = 8'h7b;
assign sbox[4] = 8'hf2;
assign sbox[5] = 8'h6b;
assign sbox[6] = 8'h6f;
assign sbox[7] = 8'hc5;
assign sbox[8] = 8'h30;
assign sbox[9] = 8'h01;
assign sbox[10] = 8'h67;
assign sbox[11] = 8'h2b;
assign sbox[12] = 8'hfe;
assign sbox[13] = 8'hd7;
assign sbox[14] = 8'hab;
assign sbox[15] = 8'h76;
assign sbox[16] = 8'hca;
assign sbox[17] = 8'h82;
assign sbox[18] = 8'hc9;
assign sbox[19] = 8'h7d;
assign sbox[20] = 8'hfa;
assign sbox[21] = 8'h59;
assign sbox[22] = 8'h47;
assign sbox[23] = 8'hf0;
assign sbox[24] = 8'had;
assign sbox[25] = 8'hd4;
assign sbox[26] = 8'ha2;
assign sbox[27] = 8'haf;
assign sbox[28] = 8'h9c;
assign sbox[29] = 8'ha4;
assign sbox[30] = 8'h72;
assign sbox[31] = 8'hc0;
assign sbox[32] = 8'hb7;
assign sbox[33] = 8'hfd;
assign sbox[34] = 8'h93;
assign sbox[35] = 8'h26;
assign sbox[36] = 8'h36;
assign sbox[37] = 8'h3f;
assign sbox[38] = 8'hf7;
assign sbox[39] = 8'hcc;
assign sbox[40] = 8'h34;
assign sbox[41] = 8'ha5;
assign sbox[42] = 8'he5;
assign sbox[43] = 8'hf1;
assign sbox[44] = 8'h71;
assign sbox[45] = 8'hd8;
assign sbox[46] = 8'h31;
assign sbox[47] = 8'h15;
assign sbox[48] = 8'h04;
assign sbox[49] = 8'hc7;
assign sbox[50] = 8'h23;
assign sbox[51] = 8'hc3;
assign sbox[52] = 8'h18;
assign sbox[53] = 8'h96;
assign sbox[54] = 8'h05;
assign sbox[55] = 8'h9a;
assign sbox[56] = 8'h07;
assign sbox[57] = 8'h12;
assign sbox[58] = 8'h80;
assign sbox[59] = 8'he2;
assign sbox[60] = 8'heb;
assign sbox[61] = 8'h27;
assign sbox[62] = 8'hb2;
assign sbox[63] = 8'h75;
assign sbox[64] = 8'h09;
assign sbox[65] = 8'h83;
assign sbox[66] = 8'h2c;
assign sbox[67] = 8'h1a;
assign sbox[68] = 8'h1b;
assign sbox[69] = 8'h6e;
assign sbox[70] = 8'h5a;
assign sbox[71] = 8'ha0;
assign sbox[72] = 8'h52;
assign sbox[73] = 8'h3b;
assign sbox[74] = 8'hd6;
assign sbox[75] = 8'hb3;
assign sbox[76] = 8'h29;
assign sbox[77] = 8'he3;
assign sbox[78] = 8'h2f;
assign sbox[79] = 8'h84;
assign sbox[80] = 8'h53;
assign sbox[81] = 8'hd1;
assign sbox[82] = 8'h00;
assign sbox[83] = 8'hed;
assign sbox[84] = 8'h20;
assign sbox[85] = 8'hfc;
assign sbox[86] = 8'hb1;
assign sbox[87] = 8'h5b;
assign sbox[88] = 8'h6a;
assign sbox[89] = 8'hcb;
assign sbox[90] = 8'hbe;
assign sbox[91] = 8'h39;
assign sbox[92] = 8'h4a;
assign sbox[93] = 8'h4c;
assign sbox[94] = 8'h58;
assign sbox[95] = 8'hcf;
assign sbox[96] = 8'hd0;
assign sbox[97] = 8'hef;
assign sbox[98] = 8'haa;
assign sbox[99] = 8'hfb;
assign sbox[100] = 8'h43;
assign sbox[101] = 8'h4d;
assign sbox[102] = 8'h33;
assign sbox[103] = 8'h85;
assign sbox[104] = 8'h45;
assign sbox[105] = 8'hf9;
assign sbox[106] = 8'h02;
assign sbox[107] = 8'h7f;
assign sbox[108] = 8'h50;
assign sbox[109] = 8'h3c;
assign sbox[110] = 8'h9f;
assign sbox[111] = 8'ha8;
assign sbox[112] = 8'h51;
assign sbox[113] = 8'ha3;
assign sbox[114] = 8'h40;
assign sbox[115] = 8'h8f;
assign sbox[116] = 8'h92;
assign sbox[117] = 8'h9d;
assign sbox[118] = 8'h38;
assign sbox[119] = 8'hf5;
assign sbox[120] = 8'hbc;
assign sbox[121] = 8'hb6;
assign sbox[122] = 8'hda;
assign sbox[123] = 8'h21;
assign sbox[124] = 8'h10;
assign sbox[125] = 8'hff;
assign sbox[126] = 8'hf3;
assign sbox[127] = 8'hd2;
assign sbox[128] = 8'hcd;
assign sbox[129] = 8'h0c;
assign sbox[130] = 8'h13;
assign sbox[131] = 8'hec;
assign sbox[132] = 8'h5f;
assign sbox[133] = 8'h97;
assign sbox[134] = 8'h44;
assign sbox[135] = 8'h17;
assign sbox[136] = 8'hc4;
assign sbox[137] = 8'ha7;
assign sbox[138] = 8'h7e;
assign sbox[139] = 8'h3d;
assign sbox[140] = 8'h64;
assign sbox[141] = 8'h5d;
assign sbox[142] = 8'h19;
assign sbox[143] = 8'h73;
assign sbox[144] = 8'h60;
assign sbox[145] = 8'h81;
assign sbox[146] = 8'h4f;
assign sbox[147] = 8'hdc;
assign sbox[148] = 8'h22;
assign sbox[149] = 8'h2a;
assign sbox[150] = 8'h90;
assign sbox[151] = 8'h88;
assign sbox[152] = 8'h46;
assign sbox[153] = 8'hee;
assign sbox[154] = 8'hb8;
assign sbox[155] = 8'h14;
assign sbox[156] = 8'hde;
assign sbox[157] = 8'h5e;
assign sbox[158] = 8'h0b;
assign sbox[159] = 8'hdb;
assign sbox[160] = 8'he0;
assign sbox[161] = 8'h32;
assign sbox[162] = 8'h3a;
assign sbox[163] = 8'h0a;
assign sbox[164] = 8'h49;
assign sbox[165] = 8'h06;
assign sbox[166] = 8'h24;
assign sbox[167] = 8'h5c;
assign sbox[168] = 8'hc2;
assign sbox[169] = 8'hd3;
assign sbox[170] = 8'hac;
assign sbox[171] = 8'h62;
assign sbox[172] = 8'h91;
assign sbox[173] = 8'h95;
assign sbox[174] = 8'he4;
assign sbox[175] = 8'h79;
assign sbox[176] = 8'he7;
assign sbox[177] = 8'hc8;
assign sbox[178] = 8'h37;
assign sbox[179] = 8'h6d;
assign sbox[180] = 8'h8d;
assign sbox[181] = 8'hd5;
assign sbox[182] = 8'h4e;
assign sbox[183] = 8'ha9;
assign sbox[184] = 8'h6c;
assign sbox[185] = 8'h56;
assign sbox[186] = 8'hf4;
assign sbox[187] = 8'hea;
assign sbox[188] = 8'h65;
assign sbox[189] = 8'h7a;
assign sbox[190] = 8'hae;
assign sbox[191] = 8'h08;
assign sbox[192] = 8'hba;
assign sbox[193] = 8'h78;
assign sbox[194] = 8'h25;
assign sbox[195] = 8'h2e;
assign sbox[196] = 8'h1c;
assign sbox[197] = 8'ha6;
assign sbox[198] = 8'hb4;
assign sbox[199] = 8'hc6;
assign sbox[200] = 8'he8;
assign sbox[201] = 8'hdd;
assign sbox[202] = 8'h74;
assign sbox[203] = 8'h1f;
assign sbox[204] = 8'h4b;
assign sbox[205] = 8'hbd;
assign sbox[206] = 8'h8b;
assign sbox[207] = 8'h8a;
assign sbox[208] = 8'h70;
assign sbox[209] = 8'h3e;
assign sbox[210] = 8'hb5;
assign sbox[211] = 8'h66;
assign sbox[212] = 8'h48;
assign sbox[213] = 8'h03;
assign sbox[214] = 8'hf6;
assign sbox[215] = 8'h0e;
assign sbox[216] = 8'h61;
assign sbox[217] = 8'h35;
assign sbox[218] = 8'h57;
assign sbox[219] = 8'hb9;
assign sbox[220] = 8'h86;
assign sbox[221] = 8'hc1;
assign sbox[222] = 8'h1d;
assign sbox[223] = 8'h9e;
assign sbox[224] = 8'he1;
assign sbox[225] = 8'hf8;
assign sbox[226] = 8'h98;
assign sbox[227] = 8'h11;
assign sbox[228] = 8'h69;
assign sbox[229] = 8'hd9;
assign sbox[230] = 8'h8e;
assign sbox[231] = 8'h94;
assign sbox[232] = 8'h9b;
assign sbox[233] = 8'h1e;
assign sbox[234] = 8'h87;
assign sbox[235] = 8'he9;
assign sbox[236] = 8'hce;
assign sbox[237] = 8'h55;
assign sbox[238] = 8'h28;
assign sbox[239] = 8'hdf;
assign sbox[240] = 8'h8c;
assign sbox[241] = 8'ha1;
assign sbox[242] = 8'h89;
assign sbox[243] = 8'h0d;
assign sbox[244] = 8'hbf;
assign sbox[245] = 8'he6;
assign sbox[246] = 8'h42;
assign sbox[247] = 8'h68;
assign sbox[248] = 8'h41;
assign sbox[249] = 8'h99;
assign sbox[250] = 8'h2d;
assign sbox[251] = 8'h0f;
assign sbox[252] = 8'hb0;
assign sbox[253] = 8'h54;
assign sbox[254] = 8'hbb;
assign sbox[255] = 8'h16;

endmodule