// this module implements a combo of sbox and tbox for a whole column
module direct_sbox_tbox(in_word, out_words);

input [0:31] in_word;
output [0:39] out_words[0:3];

wire [0:39] sbox_tbox[0:255];
wire [7:0] in_byte[0:3];
wire [0:39] mapping[0:3];

genvar i;
generate
    for(i = 0; i < 4; i++)
        begin: split_and_mapping
        // split original 32-bit column word into 4 bytes
        assign in_byte[i] = in_word[i*8:(i+1)*8-1];
        // map the "addresses" to the correct rom entry
        assign mapping[i] = sbox_tbox[in_byte[i]];
        end
endgenerate

assign out_words[0] = mapping[0];
assign out_words[1] = {mapping[1][0:7], mapping[1][8:39] >> 8 | mapping[1][8:39] << 24};
assign out_words[2] = {mapping[2][0:7], mapping[2][8:39] >> 16 | mapping[2][8:39] << 16};
assign out_words[3] = {mapping[3][0:7], mapping[3][8:39] >> 24 | mapping[3][8:39] << 8};

// hardwired implementation of the sbox_tbox mapping
assign sbox_tbox[0] = 40'h63c66363a5;
assign sbox_tbox[1] = 40'h7cf87c7c84;
assign sbox_tbox[2] = 40'h77ee777799;
assign sbox_tbox[3] = 40'h7bf67b7b8d;
assign sbox_tbox[4] = 40'hf2fff2f20d;
assign sbox_tbox[5] = 40'h6bd66b6bbd;
assign sbox_tbox[6] = 40'h6fde6f6fb1;
assign sbox_tbox[7] = 40'hc591c5c554;
assign sbox_tbox[8] = 40'h3060303050;
assign sbox_tbox[9] = 40'h0102010103;
assign sbox_tbox[10] = 40'h67ce6767a9;
assign sbox_tbox[11] = 40'h2b562b2b7d;
assign sbox_tbox[12] = 40'hfee7fefe19;
assign sbox_tbox[13] = 40'hd7b5d7d762;
assign sbox_tbox[14] = 40'hab4dababe6;
assign sbox_tbox[15] = 40'h76ec76769a;
assign sbox_tbox[16] = 40'hca8fcaca45;
assign sbox_tbox[17] = 40'h821f82829d;
assign sbox_tbox[18] = 40'hc989c9c940;
assign sbox_tbox[19] = 40'h7dfa7d7d87;
assign sbox_tbox[20] = 40'hfaeffafa15;
assign sbox_tbox[21] = 40'h59b25959eb;
assign sbox_tbox[22] = 40'h478e4747c9;
assign sbox_tbox[23] = 40'hf0fbf0f00b;
assign sbox_tbox[24] = 40'had41adadec;
assign sbox_tbox[25] = 40'hd4b3d4d467;
assign sbox_tbox[26] = 40'ha25fa2a2fd;
assign sbox_tbox[27] = 40'haf45afafea;
assign sbox_tbox[28] = 40'h9c239c9cbf;
assign sbox_tbox[29] = 40'ha453a4a4f7;
assign sbox_tbox[30] = 40'h72e4727296;
assign sbox_tbox[31] = 40'hc09bc0c05b;
assign sbox_tbox[32] = 40'hb775b7b7c2;
assign sbox_tbox[33] = 40'hfde1fdfd1c;
assign sbox_tbox[34] = 40'h933d9393ae;
assign sbox_tbox[35] = 40'h264c26266a;
assign sbox_tbox[36] = 40'h366c36365a;
assign sbox_tbox[37] = 40'h3f7e3f3f41;
assign sbox_tbox[38] = 40'hf7f5f7f702;
assign sbox_tbox[39] = 40'hcc83cccc4f;
assign sbox_tbox[40] = 40'h346834345c;
assign sbox_tbox[41] = 40'ha551a5a5f4;
assign sbox_tbox[42] = 40'he5d1e5e534;
assign sbox_tbox[43] = 40'hf1f9f1f108;
assign sbox_tbox[44] = 40'h71e2717193;
assign sbox_tbox[45] = 40'hd8abd8d873;
assign sbox_tbox[46] = 40'h3162313153;
assign sbox_tbox[47] = 40'h152a15153f;
assign sbox_tbox[48] = 40'h040804040c;
assign sbox_tbox[49] = 40'hc795c7c752;
assign sbox_tbox[50] = 40'h2346232365;
assign sbox_tbox[51] = 40'hc39dc3c35e;
assign sbox_tbox[52] = 40'h1830181828;
assign sbox_tbox[53] = 40'h96379696a1;
assign sbox_tbox[54] = 40'h050a05050f;
assign sbox_tbox[55] = 40'h9a2f9a9ab5;
assign sbox_tbox[56] = 40'h070e070709;
assign sbox_tbox[57] = 40'h1224121236;
assign sbox_tbox[58] = 40'h801b80809b;
assign sbox_tbox[59] = 40'he2dfe2e23d;
assign sbox_tbox[60] = 40'hebcdebeb26;
assign sbox_tbox[61] = 40'h274e272769;
assign sbox_tbox[62] = 40'hb27fb2b2cd;
assign sbox_tbox[63] = 40'h75ea75759f;
assign sbox_tbox[64] = 40'h091209091b;
assign sbox_tbox[65] = 40'h831d83839e;
assign sbox_tbox[66] = 40'h2c582c2c74;
assign sbox_tbox[67] = 40'h1a341a1a2e;
assign sbox_tbox[68] = 40'h1b361b1b2d;
assign sbox_tbox[69] = 40'h6edc6e6eb2;
assign sbox_tbox[70] = 40'h5ab45a5aee;
assign sbox_tbox[71] = 40'ha05ba0a0fb;
assign sbox_tbox[72] = 40'h52a45252f6;
assign sbox_tbox[73] = 40'h3b763b3b4d;
assign sbox_tbox[74] = 40'hd6b7d6d661;
assign sbox_tbox[75] = 40'hb37db3b3ce;
assign sbox_tbox[76] = 40'h295229297b;
assign sbox_tbox[77] = 40'he3dde3e33e;
assign sbox_tbox[78] = 40'h2f5e2f2f71;
assign sbox_tbox[79] = 40'h8413848497;
assign sbox_tbox[80] = 40'h53a65353f5;
assign sbox_tbox[81] = 40'hd1b9d1d168;
assign sbox_tbox[82] = 40'h0000000000;
assign sbox_tbox[83] = 40'hedc1eded2c;
assign sbox_tbox[84] = 40'h2040202060;
assign sbox_tbox[85] = 40'hfce3fcfc1f;
assign sbox_tbox[86] = 40'hb179b1b1c8;
assign sbox_tbox[87] = 40'h5bb65b5bed;
assign sbox_tbox[88] = 40'h6ad46a6abe;
assign sbox_tbox[89] = 40'hcb8dcbcb46;
assign sbox_tbox[90] = 40'hbe67bebed9;
assign sbox_tbox[91] = 40'h397239394b;
assign sbox_tbox[92] = 40'h4a944a4ade;
assign sbox_tbox[93] = 40'h4c984c4cd4;
assign sbox_tbox[94] = 40'h58b05858e8;
assign sbox_tbox[95] = 40'hcf85cfcf4a;
assign sbox_tbox[96] = 40'hd0bbd0d06b;
assign sbox_tbox[97] = 40'hefc5efef2a;
assign sbox_tbox[98] = 40'haa4faaaae5;
assign sbox_tbox[99] = 40'hfbedfbfb16;
assign sbox_tbox[100] = 40'h43864343c5;
assign sbox_tbox[101] = 40'h4d9a4d4dd7;
assign sbox_tbox[102] = 40'h3366333355;
assign sbox_tbox[103] = 40'h8511858594;
assign sbox_tbox[104] = 40'h458a4545cf;
assign sbox_tbox[105] = 40'hf9e9f9f910;
assign sbox_tbox[106] = 40'h0204020206;
assign sbox_tbox[107] = 40'h7ffe7f7f81;
assign sbox_tbox[108] = 40'h50a05050f0;
assign sbox_tbox[109] = 40'h3c783c3c44;
assign sbox_tbox[110] = 40'h9f259f9fba;
assign sbox_tbox[111] = 40'ha84ba8a8e3;
assign sbox_tbox[112] = 40'h51a25151f3;
assign sbox_tbox[113] = 40'ha35da3a3fe;
assign sbox_tbox[114] = 40'h40804040c0;
assign sbox_tbox[115] = 40'h8f058f8f8a;
assign sbox_tbox[116] = 40'h923f9292ad;
assign sbox_tbox[117] = 40'h9d219d9dbc;
assign sbox_tbox[118] = 40'h3870383848;
assign sbox_tbox[119] = 40'hf5f1f5f504;
assign sbox_tbox[120] = 40'hbc63bcbcdf;
assign sbox_tbox[121] = 40'hb677b6b6c1;
assign sbox_tbox[122] = 40'hdaafdada75;
assign sbox_tbox[123] = 40'h2142212163;
assign sbox_tbox[124] = 40'h1020101030;
assign sbox_tbox[125] = 40'hffe5ffff1a;
assign sbox_tbox[126] = 40'hf3fdf3f30e;
assign sbox_tbox[127] = 40'hd2bfd2d26d;
assign sbox_tbox[128] = 40'hcd81cdcd4c;
assign sbox_tbox[129] = 40'h0c180c0c14;
assign sbox_tbox[130] = 40'h1326131335;
assign sbox_tbox[131] = 40'hecc3ecec2f;
assign sbox_tbox[132] = 40'h5fbe5f5fe1;
assign sbox_tbox[133] = 40'h97359797a2;
assign sbox_tbox[134] = 40'h44884444cc;
assign sbox_tbox[135] = 40'h172e171739;
assign sbox_tbox[136] = 40'hc493c4c457;
assign sbox_tbox[137] = 40'ha755a7a7f2;
assign sbox_tbox[138] = 40'h7efc7e7e82;
assign sbox_tbox[139] = 40'h3d7a3d3d47;
assign sbox_tbox[140] = 40'h64c86464ac;
assign sbox_tbox[141] = 40'h5dba5d5de7;
assign sbox_tbox[142] = 40'h193219192b;
assign sbox_tbox[143] = 40'h73e6737395;
assign sbox_tbox[144] = 40'h60c06060a0;
assign sbox_tbox[145] = 40'h8119818198;
assign sbox_tbox[146] = 40'h4f9e4f4fd1;
assign sbox_tbox[147] = 40'hdca3dcdc7f;
assign sbox_tbox[148] = 40'h2244222266;
assign sbox_tbox[149] = 40'h2a542a2a7e;
assign sbox_tbox[150] = 40'h903b9090ab;
assign sbox_tbox[151] = 40'h880b888883;
assign sbox_tbox[152] = 40'h468c4646ca;
assign sbox_tbox[153] = 40'heec7eeee29;
assign sbox_tbox[154] = 40'hb86bb8b8d3;
assign sbox_tbox[155] = 40'h142814143c;
assign sbox_tbox[156] = 40'hdea7dede79;
assign sbox_tbox[157] = 40'h5ebc5e5ee2;
assign sbox_tbox[158] = 40'h0b160b0b1d;
assign sbox_tbox[159] = 40'hdbaddbdb76;
assign sbox_tbox[160] = 40'he0dbe0e03b;
assign sbox_tbox[161] = 40'h3264323256;
assign sbox_tbox[162] = 40'h3a743a3a4e;
assign sbox_tbox[163] = 40'h0a140a0a1e;
assign sbox_tbox[164] = 40'h49924949db;
assign sbox_tbox[165] = 40'h060c06060a;
assign sbox_tbox[166] = 40'h244824246c;
assign sbox_tbox[167] = 40'h5cb85c5ce4;
assign sbox_tbox[168] = 40'hc29fc2c25d;
assign sbox_tbox[169] = 40'hd3bdd3d36e;
assign sbox_tbox[170] = 40'hac43acacef;
assign sbox_tbox[171] = 40'h62c46262a6;
assign sbox_tbox[172] = 40'h91399191a8;
assign sbox_tbox[173] = 40'h95319595a4;
assign sbox_tbox[174] = 40'he4d3e4e437;
assign sbox_tbox[175] = 40'h79f279798b;
assign sbox_tbox[176] = 40'he7d5e7e732;
assign sbox_tbox[177] = 40'hc88bc8c843;
assign sbox_tbox[178] = 40'h376e373759;
assign sbox_tbox[179] = 40'h6dda6d6db7;
assign sbox_tbox[180] = 40'h8d018d8d8c;
assign sbox_tbox[181] = 40'hd5b1d5d564;
assign sbox_tbox[182] = 40'h4e9c4e4ed2;
assign sbox_tbox[183] = 40'ha949a9a9e0;
assign sbox_tbox[184] = 40'h6cd86c6cb4;
assign sbox_tbox[185] = 40'h56ac5656fa;
assign sbox_tbox[186] = 40'hf4f3f4f407;
assign sbox_tbox[187] = 40'heacfeaea25;
assign sbox_tbox[188] = 40'h65ca6565af;
assign sbox_tbox[189] = 40'h7af47a7a8e;
assign sbox_tbox[190] = 40'hae47aeaee9;
assign sbox_tbox[191] = 40'h0810080818;
assign sbox_tbox[192] = 40'hba6fbabad5;
assign sbox_tbox[193] = 40'h78f0787888;
assign sbox_tbox[194] = 40'h254a25256f;
assign sbox_tbox[195] = 40'h2e5c2e2e72;
assign sbox_tbox[196] = 40'h1c381c1c24;
assign sbox_tbox[197] = 40'ha657a6a6f1;
assign sbox_tbox[198] = 40'hb473b4b4c7;
assign sbox_tbox[199] = 40'hc697c6c651;
assign sbox_tbox[200] = 40'he8cbe8e823;
assign sbox_tbox[201] = 40'hdda1dddd7c;
assign sbox_tbox[202] = 40'h74e874749c;
assign sbox_tbox[203] = 40'h1f3e1f1f21;
assign sbox_tbox[204] = 40'h4b964b4bdd;
assign sbox_tbox[205] = 40'hbd61bdbddc;
assign sbox_tbox[206] = 40'h8b0d8b8b86;
assign sbox_tbox[207] = 40'h8a0f8a8a85;
assign sbox_tbox[208] = 40'h70e0707090;
assign sbox_tbox[209] = 40'h3e7c3e3e42;
assign sbox_tbox[210] = 40'hb571b5b5c4;
assign sbox_tbox[211] = 40'h66cc6666aa;
assign sbox_tbox[212] = 40'h48904848d8;
assign sbox_tbox[213] = 40'h0306030305;
assign sbox_tbox[214] = 40'hf6f7f6f601;
assign sbox_tbox[215] = 40'h0e1c0e0e12;
assign sbox_tbox[216] = 40'h61c26161a3;
assign sbox_tbox[217] = 40'h356a35355f;
assign sbox_tbox[218] = 40'h57ae5757f9;
assign sbox_tbox[219] = 40'hb969b9b9d0;
assign sbox_tbox[220] = 40'h8617868691;
assign sbox_tbox[221] = 40'hc199c1c158;
assign sbox_tbox[222] = 40'h1d3a1d1d27;
assign sbox_tbox[223] = 40'h9e279e9eb9;
assign sbox_tbox[224] = 40'he1d9e1e138;
assign sbox_tbox[225] = 40'hf8ebf8f813;
assign sbox_tbox[226] = 40'h982b9898b3;
assign sbox_tbox[227] = 40'h1122111133;
assign sbox_tbox[228] = 40'h69d26969bb;
assign sbox_tbox[229] = 40'hd9a9d9d970;
assign sbox_tbox[230] = 40'h8e078e8e89;
assign sbox_tbox[231] = 40'h94339494a7;
assign sbox_tbox[232] = 40'h9b2d9b9bb6;
assign sbox_tbox[233] = 40'h1e3c1e1e22;
assign sbox_tbox[234] = 40'h8715878792;
assign sbox_tbox[235] = 40'he9c9e9e920;
assign sbox_tbox[236] = 40'hce87cece49;
assign sbox_tbox[237] = 40'h55aa5555ff;
assign sbox_tbox[238] = 40'h2850282878;
assign sbox_tbox[239] = 40'hdfa5dfdf7a;
assign sbox_tbox[240] = 40'h8c038c8c8f;
assign sbox_tbox[241] = 40'ha159a1a1f8;
assign sbox_tbox[242] = 40'h8909898980;
assign sbox_tbox[243] = 40'h0d1a0d0d17;
assign sbox_tbox[244] = 40'hbf65bfbfda;
assign sbox_tbox[245] = 40'he6d7e6e631;
assign sbox_tbox[246] = 40'h42844242c6;
assign sbox_tbox[247] = 40'h68d06868b8;
assign sbox_tbox[248] = 40'h41824141c3;
assign sbox_tbox[249] = 40'h99299999b0;
assign sbox_tbox[250] = 40'h2d5a2d2d77;
assign sbox_tbox[251] = 40'h0f1e0f0f11;
assign sbox_tbox[252] = 40'hb07bb0b0cb;
assign sbox_tbox[253] = 40'h54a85454fc;
assign sbox_tbox[254] = 40'hbb6dbbbbd6;
assign sbox_tbox[255] = 40'h162c16163a;

endmodule